package simple_req_ack_uvc_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"

`include "simple_req_ack_transaction.sv"
`include "simple_req_ack_uvc_cfg.sv"
`include "simple_req_ack_monitor.sv"
`include "simple_req_ack_sequencer.sv"
`include "simple_req_ack_driver.sv"
`include "simple_req_ack_agent.sv"
`include "simple_req_ack_seq_lib.sv"


endpackage: simple_req_ack_uvc_pkg

